module decodetest;
